module test(in,led);
input in;
output led;
	assign led = in;
endmodule
