`timescale 1ns / 1ps

module test(in,led);
assign led = in;
endmodule
